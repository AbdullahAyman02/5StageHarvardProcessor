LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY EPC_TB IS
END ENTITY;

ARCHITECTURE EPC_TB_ARCH OF EPC_TB IS
    COMPONENT EPC
        PORT(
            OVERFLOW_PC  : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            PROTECTED_PC : IN STD_LOGIC_VECTOR(31 DOWNTO 0);

            OVERFLOW_FLAG : IN STD_LOGIC;
            PROTECTED_FLAG  : IN STD_LOGIC;

            EPC_PC : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
            EPC_FLAG : OUT STD_LOGIC
        );
    END COMPONENT;

    SIGNAL OVERFLOW_PC  : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL PROTECTED_PC : STD_LOGIC_VECTOR(31 DOWNTO 0);

    SIGNAL OVERFLOW_FLAG : STD_LOGIC;
    SIGNAL PROTECTED_FLAG  : STD_LOGIC;

    SIGNAL EPC_PC : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL EPC_FLAG : STD_LOGIC;

BEGIN
    UUT: EPC PORT MAP(
        OVERFLOW_PC => OVERFLOW_PC,
        PROTECTED_PC => PROTECTED_PC,
        OVERFLOW_FLAG => OVERFLOW_FLAG,
        PROTECTED_FLAG => PROTECTED_FLAG,
        EPC_PC => EPC_PC,
        EPC_FLAG => EPC_FLAG
    );

    TEST: PROCESS
    BEGIN
        -- '1' OVERFLOW, '0' PROTECTED
        
        OVERFLOW_PC <= X"00000001";
        PROTECTED_PC <= X"00000002";
        
        -- TEST CASE 1: OVERFLOW_FLAG = '0', PROTECTED_FLAG = '0'
        OVERFLOW_FLAG <= '0';
        PROTECTED_FLAG <= '0';
        WAIT FOR 10 ns;
        ASSERT (EPC_PC = X"00000002" AND EPC_FLAG = '0') REPORT "TEST CASE 1 FAILED" SEVERITY ERROR;

        -- TEST CASE 2: OVERFLOW_FLAG = '0', PROTECTED_FLAG = '1'
        OVERFLOW_FLAG <= '0';
        PROTECTED_FLAG <= '1';
        WAIT FOR 10 ns;
        ASSERT (EPC_PC = X"00000002" AND EPC_FLAG = '0') REPORT "TEST CASE 2 FAILED" SEVERITY ERROR;

        -- TEST CASE 3: OVERFLOW_FLAG = '1', PROTECTED_FLAG = '0'
        OVERFLOW_FLAG <= '1';
        PROTECTED_FLAG <= '0';
        WAIT FOR 10 ns;
        ASSERT (EPC_PC = X"00000001" AND EPC_FLAG = '1') REPORT "TEST CASE 3 FAILED" SEVERITY ERROR;

        -- TEST CASE 4: OVERFLOW_FLAG = '1', PROTECTED_FLAG = '1'
        OVERFLOW_FLAG <= '1';
        PROTECTED_FLAG <= '1';
        WAIT FOR 10 ns;
        ASSERT (EPC_PC = X"00000002" AND EPC_FLAG = '0') REPORT "TEST CASE 4 FAILED" SEVERITY ERROR;

        WAIT;
    END PROCESS TEST;
END ARCHITECTURE EPC_TB_ARCH;